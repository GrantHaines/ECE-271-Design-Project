/*

	Top-level module for the design project

*/

module top-level();



endmodule