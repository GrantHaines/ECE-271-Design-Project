module comp(input logic [5:0] a, b,
            output logic gt);
 
   assign gt = (a > b);

endmodule 